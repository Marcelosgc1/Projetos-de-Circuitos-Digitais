module decoder_irrigation(
input Bit0,
input Bit1,
output a,
output b,
output c,
output d,
output e,
output f,
output g,
output digit
);

	
	//01 -> A, B, C, E, F, G
	//10 -> A, C, D, E, F
	//11 -> A, B, C, D, E, F
	
	
	
	
	
	
	
endmodule 
