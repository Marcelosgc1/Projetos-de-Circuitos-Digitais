module timer();

endmodule
