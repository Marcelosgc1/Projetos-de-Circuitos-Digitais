module stopwatch();

endmodule
